----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/15/2018 05:51:44 PM
-- Design Name: 
-- Module Name: InstructionMemory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity InstructionMemory is

PORT ( A: in STD_LOGIC_VECTOR(31 DOWNTO 0);
 	   RD: out STD_LOGIC_VECTOR(31 DOWNTO 0));

end InstructionMemory;

architecture Behavioral of InstructionMemory is

TYPE rom IS ARRAY (0 TO 683) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
CONSTANT imem: 
rom:=rom'(  

--------------- skey generation --------------------------------

"00000000","00000000","00000000","00000011",       -- SUB R0,R0,R0            -- INSTR1  --
"00000000","00100001","00001000","00000011",       -- SUB R1,R1,R1            -- INSTR2  -- K_CNT = 0
"00000000","01000010","00010000","00000011",       -- SUB R2,R2,R2            -- INSTR3  -- I_CNT = 0
"00000000","01100011","00011000","00000011",       -- SUB R3,R3,R3            -- INSTR4  -- J_CNT = 0
"00000001","01101011","01011000","00000011",       -- SUB R11,R11,R11         -- INSTR5  -- NUMBER OF TIMES ROTATION IS CALLED

"00011100","00000100","00000000","01110100",       -- LB R0,R4,x"0074"        -- INSTR6  -- R4 = A
"00011100","00000101","00000000","01111000",       -- LB R0,R5,x"0078"        -- INSTR7  -- R5 = B
"00011100","00001100","00000000","01110000",       -- LB R0,R12,x"0070"       -- INSTR8  -- R12 = x"80000000"

"00000000","01000010","01101000","00000001",	   --ADD R2,R2,R13            -- INSTR9  -- R13 = 2i
"00000001","10101101","01101000","00000001",	   --ADD R13,R13,R13          -- INSTR10  -- R13 = 4i
"00011101","10100110","00000000","01111100",       -- LB R13,R6,x"007C"       -- INSTR11 -- R6 = s[i]
"00000000","01100011","01110000","00000001",	   --ADD R3,R3,R14            -- INSTR12  -- R14 = 2j
"00000001","11001110","01110000","00000001",	   --ADD R14,R14,R14          -- INSTR13  -- R14 = 4j
"00011101","11000111","00000000","11100100",       -- LB R14,R7,x"00E4"       -- INSTR14 -- R7 = L[j]

"00000000","10000101","01000000","00000001",       -- ADD R4,R5,R8            -- INSTR15 -- R8 = A+B
"00000001","00000110","01111000","00000001",       -- ADD R8,R6,R15           -- INSTR16 -- R15 = s[i]+A+B
"00000100","00001000","00000000","00000011",       -- ADDI R0,R8,x"0003"      -- INSTR17 -- R8 = 3
"00110000","00000000","00000000","00101101",       -- JMP (INSTR = 46)        -- INSTR18 -- JUMP TO skey_ROTATION 
"00101000","00010000","00000000","00000110",       -- BEQ R0,R16,(INSTR = 26) -- INSTR19 -- UPDATING A/B IN THE ITERATION
"00000000","00001111","00110000","00000001",       -- ADD R0,R15,R6           -- INSTR20 -- s[i] = (s[i]+A+B)<<<3
"00100001","10100110","00000000","01111100",       -- SB R13,R6,x"007C"       -- INSTR21 -- STORE IN s[i]
"00000000","00001111","00100000","00000001",       -- ADD R0,R15,R4           -- INSTR22 -- A = (s[i]+A+B)<<<3
"00000000","10000101","01000000","00000001",       -- ADD R4,R5,R8            -- INSTR23 -- R8 = A+B
"00000001","00000111","01111000","00000001",       -- ADD R8,R7,R15           -- INSTR24 -- R15 = L[j]+A+B
"00110000","00000000","00000000","00101101",       -- JMP (INSTR = 46)        -- INSTR25 -- JUMP TO ROTATION 
"00000000","00001111","00111000","00000001",       -- ADD R0,R15,R7           -- INSTR26 -- L[j] = (L[j]+A+B)<<<(A+B)
"00100001","11000111","00000000","11100100",       -- SB R14,R7,x"00E4"       -- INSTR27 -- STORE IN L[j]
"00000000","00001111","00101000","00000001",       -- ADD R0,R15,R5           -- INSTR28 -- B = (L[j]+A+B)<<<(A+B)

"00000100","00001010","00000000","01001101",       -- ADDI R0,R10,x"004D"     -- INSTR29 -- R10 = 77  
"00101000","00101010","00000000","00001100",       -- BEQ R1,R10,(INSTR = 43) -- INSTR30 -- JUMP TO HALT
"00000100","00100001","00000000","00000001",       -- ADDI R1,R1,x"0001"      -- INSTR31 -- K_CNT = K_CNT +1

"00000100","00001010","00000000","00011001",       -- ADDI R0,R10,x"0019"     -- INSTR32 -- R10 = 25  
"00101100","01001010","00000000","00000010",       -- BNEQ R2,R10,(INSTR = 36)-- INSTR33 -- 
"00000000","01000010","00010000","00000011",       -- SUB R2,R2,R2            -- INSTR34 -- I_CNT = 0
"00110000","00000000","00000000","00100100",       -- JMP (INSTR = 37)        -- INSTR35 -- 
"00000100","01000010","00000000","00000001",       -- ADDI R2,R2,x"0001"      -- INSTR36 -- I_CNT = I_CNT +1

"00000100","00001010","00000000","00000011",       -- ADDI R0,R10,x"0003"     -- INSTR37 -- R10 = 3  
"00101100","01101010","00000000","00000010",       -- BNEQ R3,R10,(INSTR = 41)-- INSTR38 -- 
"00000000","01100011","00011000","00000011",       -- SUB R3,R3,R3            -- INSTR39 -- J_CNT = 0
"00110000","00000000","00000000","00001000",       -- JMP (INSTR = 9)         -- INSTR40 -- 
"00000100","01100011","00000000","00000001",       -- ADDI R3,R3,x"0001"      -- INSTR41 -- J_CNT = J_CNT +1

"00110000","00000000","00000000","00001000",       -- JMP (INSTR = 9)         -- INSTR42-- 
"00011100","00010100","00000001","00000100",       -- LB R0,R20,x"0104"        -- INSTR43  -- R4 = E/D
"00101000","00010100","00000000","01001001",       -- BEQ R0,R20,(INSTR = 118) -- INSTR44 -- JUMP TO ENCRYPTION
"00110000","00000000","00000000","00111111",       -- JMP (INSTR = 64))       -- INSTR45 -- JMP to DECRYPTion
-------------------skey_ROTATION-------------------------

"00000100","00010000","00000000","00011111",	--ADDI R0,R16, x"001F"    -- INSTR 46 -- 
"00000001","00010000","10001000","00000101",	--AND R8,R16,R17          -- INSTR 47 -- LAST 5 BITS OF R7
"00000110","00010000","00000000","00000001",	--ADDI R16,R16, x"0001"   -- INSTR 48 -- R16 = 32 IN DECIMAL
"00000010","00010001","10001000","00000011",	--SUB R16,R17,R17         -- INSTR 49 -- R17 = 32 - LAST 5 BITS OF R7 
"00000010","01110011","10011000","00000011",	--SUB R19,R19,R19         -- INSTR 50 -- ROTATION COUNTER
"00000100","00010000","00000000","00000001",	--ADDI R0,R16, x"0001"    -- INSTR 51 -- 
"00000001","11110000","10010000","00000101",	--AND R15,R16,R18         -- INSTR 52 -- CHECK THE LAST BIT OF R15
"00000110","01110011","00000000","00000001",	--ADDI R19,R19, x"0001"   -- INSTR 53 -- INCREMENT ROTATION COUNTER
"00010101","11101111","00000000","00000001",	--SHR R15,R15, x"0001"    -- INSTR 54 -- SHIFT RIGHT BY ONE BIT
"00101010","01010000","00000000","00000010",	--BEQ R18,R16,(INSTR = 58)-- INSTR 55 -- IF THE LAST BIT IS 1, BRANCH TO ADDING 1 IN THE MSB
"00101010","01110001","00000000","00000100",	--BEQ R19,R17,(INSTR = 61)-- INSTR 56 -- END OF ROTATION CHECK
"00110000","00000000","00000000","00110011",	--JMP (INSTR = 52)        -- INSTR 57 -- NEXT Last bit and then SHR 
"00000001","11101100","01111000","00000001",	--ADD R15,R12,R15         -- INSTR 58 -- ADD x"80000000" TO R15
"00101010","01110001","00000000","00000001",	--BEQ R19,R17,(INSTR = 61)-- INSTR 59 -- END OF ROTATION CHECK
"00110000","00000000","00000000","00110011",	--JMP (INSTR = 52)        -- INSTR 60 -- NEXT SHR
"00000101","01101011","00000000","00000001",	--ADDI R11,R11, x"0001"   -- INSTR 61 -- NUMBER OF TIMES ROTATION IS CALLED
"00000001","01110000","10000000","00000101",	--AND R11,R16,R16         -- INSTR 62 -- LAST BIT OF R4
"00110000","00000000","00000000","00010010",    --JMP (INSTR = 19)        -- INSTR 63 -- JUMP BACK TO MAIN ROUTINE 

--------------------Decryption -------------------
"00000000","00000000","00000000","00000011",	--SUB R0,R0,R0            -- INSTR 64 -- R0 = 0
"00011100","00000001","00000000","00000100",	--LB R0,R1, x"0004"       -- INSTR 65 -- B_in
"00011100","00000010","00000000","00000000",	--LB R0,R2, x"0000"       -- INSTR 66 -- A_in
"00011100","00000110","00000000","01110000",	--LB R0,R6, x"0070 "      -- INSTR 67 -- R6 = x"80000000"
"00000001","00001000","01000000","00000011",	--SUB R8,R8,R8            -- INSTR 68 -- R8 = 0
"00000100","00000011","00000000","00001100",	--ADDI R0,R3,x"000C"      -- INSTR 69 -- R3 = 12, RC5 LOOP COUNTER 
"00000000","01100011","00100000","00000001",	--ADD R3,R3,R4            -- INSTR 70 -- R4 = 2i
"00000000","10000100","00100000","00000001",	--ADD R4,R4,R4            -- INSTR 71 -- R4 = 4i
"00000000","10000100","00100000","00000001",	--ADD R4,R4,R4            -- INSTR 72 -- R4 = 8i	
"00011100","10000101","00000000","10000000",	--LB R4,R5, x"0080"       -- INSTR 73 -- s[2i+1]
"00000000","00100101","00001000","00000011",	--SUB R1,R5,R1            -- INSTR 74 -- B = B - s[2i+1]
"00000000","00000001","01111000","00000001",	--ADD R0,R1,R15           -- INSTR 75 -- FIRST INPUT FOR ROTATION SUBROUTINE
"00000000","00000010","00111000","00000001",	--ADD R0,R2,R7            -- INSTR 76 -- SECOND INPUT FOR ROTATION SUBROUTINE
"00110000","00000000","00000000","01011111",	--JMP (INSTR = 96)        -- INSTR 77 -- JUMP TO ROTATION
"00101000","00010000","00000000","00000110",	--BEQ R0,R16,(INSTR = 85) -- INSTR 78 -- UPDATING A/B INSIDE THE ITERATION
"00000000","00001111","00001000","00000001",	--ADD R0,R15,R1           -- INSTR 79 -- B = ((B-s[2i+1])>>A) XOR A
"00011100","10000101","00000000","01111100",	--LB R4,R5, x"007C"       -- INSTR 80 -- s[2i]
"00000000","01000101","00010000","00000011",	--SUB R2,R5,R2            -- INSTR 81 -- A = A - s[2i]
"00000000","00000010","01111000","00000001",	--ADD R0,R2,R15           -- INSTR 82 -- FIRST INPUT FOR ROTATION SUBROUTINE
"00000000","00000001","00111000","00000001",	--ADD R0,R1,R7            -- INSTR 83 -- SECOND INPUT FOR ROTATION SUBROUTINE
"00110000","00000000","00000000","01011111",	--JMP (INSTR = 96)        -- INSTR 84 -- JUMP TO ROTATION
"00000000","00001111","00010000","00000001",	--ADD R0,R15,R2           -- INSTR 85 -- A = ((A-s[2i])>>B) XOR B
"00001000","01100011","00000000","00000001",	--SUBI R3,R3,x"0001"      -- INSTR 86 -- RC5 LOOP COUNTER DECREMENTATION
"00101000","00000011","00000000","00000001",	--BEQ R0,R3,(INSTR = 89)  -- INSTR 87 -- END OF RC5 LOOP 
"00110000","00000000","00000000","01000101",	--JMP (INSTR = 70)        -- INSTR 88 -- JUMP TO NEXT ITERATION
"00011100","00001001","00000000","01111100",	--LB R0,R9,x"007C"        -- INSTR 89 -- s[0]
"00011100","00001010","00000000","10000000",	--LB R0,R10,x"0080"       -- INSTR 90 -- s[1]
"00000000","00101010","00001000","00000011",	--SUB R1,R10,R1           -- INSTR 91 -- B = B - s[1]
"00000000","01001001","00010000","00000011",	--SUB R2,R9,R2            -- INSTR 92 -- A = A - s[0]
"00100000","00000001","00000000","11110100",    --SB R0,R1,x"00f4"        -- INSTR 93
"00100000","00000010","00000000","11111000",    --SB R0,R2,x"00f8"        -- INSTR 94
"11111100","00000000","00000000","00000000",	--HALT                    -- INSTR 95 -- Halt
		
-------------------- ROTATION -----------------
				
"00000100","00010000","00000000","00011111",	--ADDI R0,R16, x"001F"     -- INSTR 96 -- 
"00000000","11110000","10001000","00000101",	--AND R7,R16,R17           -- INSTR 97 -- LAST 5 BITS OF R7
"00000010","01010010","10010000","00000011",	--SUB R18,R18,R18          -- INSTR 98 -- ROTATION COUNTER
"00000100","00010000","00000000","00000001",	--ADDI R0,R16, x"0001"     -- INSTR 99 -- 	
"00101010","01010001","00000000","00001001",	--BEQ R18,R17,(INSTR = 110)-- INSTR 100 -- END OF ROTATION CHECK if last 5 bits are 0			
"00000001","11110000","10011000","00000101",	--AND R15,R16,R19          -- INSTR 101 -- CHECK THE LAST BIT OF R15
"00000110","01010010","00000000","00000001",	--ADDI R18,R18, x"0001"    -- INSTR 102 -- INCREMENT ROTATION COUNTER
"00010101","11101111","00000000","00000001",	--SHR R15,R15, x"0001"     -- INSTR 103 -- SHIFT RIGHT BY ONE BIT
"00101010","01110000","00000000","00000010",	--BEQ R19,R16,(INSTR = 107)-- INSTR 104 -- IF THE LAST BIT IS 1, BRANCH TO ADDING 1 IN THE MSB
"00101010","01010001","00000000","00000100",	--BEQ R18,R17,(INSTR = 110)-- INSTR 105 -- END OF ROTATION CHECK
"00110000","00000000","00000000","01100100",	--JMP (INSTR = 101)        -- INSTR 106 -- NEXT SHR 
"00000001","11100110","01111000","00000001",	--ADD R15,R6,R15           -- INSTR 107 -- ADD x"80000000" TO R15
"00101010","01010001","00000000","00000001",	--BEQ R18,R17,(INSTR = 110)-- INSTR 108 -- END OF ROTATION CHECK
"00110000","00000000","00000000","01100100",	--JMP (INSTR = 101)        -- INSTR 109 -- NEXT SHR 

-------------------- XOR -------------------

"00000001","11101111","01011000","00001001",	--NOR R15,R15,R11          -- INSTR 110 -- R15_BAR
"00000000","11100111","01100000","00001001",	--NOR R7,R7,R12            -- INSTR 111 -- R7_BAR
"00000001","11101100","01101000","00000101",	--AND R15,R12,R13          -- INSTR 112 -- R15.R7_BAR
"00000000","11101011","01110000","00000101",	--AND R7,R11,R14           -- INSTR 113 -- R7.R15_BAR 
"00000001","10101110","01111000","00000111",	--OR R13,R14,R15           -- INSTR 114 -- XOR
"00000101","00001000","00000000","00000001",	--ADDI R8,R8,x"0001"       -- INSTR 115 -- NUMBER OF TIMES XOR IS CALLED
"00000001","00010000","10000000","00000101",	--AND R8,R16,R16           -- INSTR 116 -- LAST BIT OF R8
"00110000","00000000","00000000","01001101",	--JMP (INSTR = 78)         -- INSTR 117 -- JUMP BACK TO MAIN ROUTINE


---------------------ENCRYPTION---------------------------------

"00000000","00000000","00000000","00000011",	--SUB R0,R0,R0            -- INSTR 118  -- R0 = 0
"00011100","00000001","00000000","00000000",	--LB R0,R1, x"0000"       -- INSTR 119  -- A_in
"00011100","00000010","00000000","00000100",	--LB R0,R2, x"0004"       -- INSTR 120  -- B_in
"00011100","00000011","00000000","01111100",    --LB R0,R3, x"007C"       -- INSTR 121  -- s[0]
"00011100","00000100","00000000","10000000",	--LB R0,R4, x"0080"       -- INSTR 122  -- s[1]
"00000000","00100011","00101000","00000001",	--ADD R1,R3,R5            -- INSTR 123 -- A = A_in + s[0]
"00000000","01000100","00110000","00000001",	--ADD R2,R4,R6            -- INSTR 124 -- B = B_in + s[1]
"00011100","00000011","00000000","01110000",	--LB R0,R3, x"0070"       -- INSTR 125 -- R3 = x"80000000" FOR ROTATION
"00000000","00100001","00001000","00000011",	--SUB R1,R1,R1            -- INSTR 126 -- R1 = 0 
"00000000","10000100","00100000","00000011",	--SUB R4,R4,R4            -- INSTR 127 -- R4 = 0
"00000100","00000010","00000000","00001100",	--ADDI R0,R2, x"000C"     -- INSTR 128 -- R2 = 12, RC5 LOOP COUNTER CHECK
"00000100","00100001","00000000","00000001",	--ADDI R1,R1, x"0001"     -- INSTR 129 -- R1 = R1+1, RC5 LOOP COUNTER 
"00000000","00100001","01001000","00000001",	--ADD R1,R1,R9            -- INSTR 130 -- R9 = 2i
"00000001","00101001","01001000","00000001",	--ADD R9,R9,R9            -- INSTR 131 -- R9 = 4i
"00000001","00101001","01001000","00000001",	--ADD R9,R9,R9            -- INSTR 132 -- R9 = 8i
"00000000","00000110","00111000","00000001",	--ADD R0,R6,R7            -- INSTR 133 -- SECOND INPUT FOR XOR SUBROUTINE
"00110000","00000000","00000000","10010100",	--JMP (INSTR = 149)       -- INSTR 134 -- JUMP TO XOR 
"00101000","00010000","00000000","00000110",	--BEQ R0,R16,(INSTR = 142)-- INSTR 135 -- UPDATING A/B INSIDE THE ITERATION
"00011101","00101010","00000000","01111100",	--LB R9,R10, x"007C"      -- INSTR 136 -- s[2i]
"00000001","11101010","00101000","00000001",	--ADD R15,R10,R5          -- INSTR 137 -- A = A_ROT + s[2i]
"00100000","00000101","00000001","00000000",    --SB R0,R5,x"0100"       -- INSTR 138
"00100000","00000101","00000000","00000000",    --SB R0,R5,x"0000"       -- INSTR 139
"00000000","00000101","00111000","00000001",	--ADD R0,R5,R7            -- INSTR 140 -- SECOND INPUT FOR XOR SUBROUTINE
"00110000","00000000","00000000","10010100",	--JMP (INSTR = 149)       -- INSTR 141 -- JUMP TO XOR
"00011101","00101010","00000000","10000000",	--LB R9,R10, x"0080"      -- INSTR 142 -- s[2i+1]
"00000001","11101010","00110000","00000001",	--ADD R15,R10,R6          -- INSTR 143 -- B = B_ROT + s[2i+1]
"00100000","00000110","00000000","11111100",    --SB R0,R6,x"00FC"       -- INSTR 144 
"00100000","00000110","00000000","00000100",    --SB R0,R6,x"0004"       -- INSTR 145 
"00101000","00100010","00000000","00000001",	--BEQ R1,R2,(INSTR = 148) -- INSTR 146 -- END OF RC5 LOOP (HALT)
"00110000","00000000","00000000","10000000",	--JMP (INSTR = 129)       -- INSTR 147 -- JUMP TO RC5 LOOP COUNTER INCREMENTATION
"00110000","00000000","00000000","00111111",	--JMP (INSTR = 64)        -- INSTR 148 -- JUMP TO Decryption
                                                                                   
-----------------------XOR----------------------------------------                                      
                                                                                   
"00000000","10100101","01011000","00001001",	--NOR R5,R5,R11           -- INSTR 149        -- R5_BAR
"00000000","11000110","01100000","00001001",	--NOR R6,R6,R12           -- INSTR 150       -- R6_BAR
"00000000","10101100","01101000","00000101",	--AND R5,R12,R13          -- INSTR 151       -- R5.R6_BAR
"00000000","11001011","01110000","00000101",	--AND R6,R11,R14          -- INSTR 152 -- -- R6.R5_BAR 
"00000001","10101110","01111000","00000111",	--OR R13,R14,R15          -- INSTR 153 -- -- XOR
                                                                                    
-----------------------ROTATION-----------------------------------                                       
                                                                                    
"00000100","00010000","00000000","00011111",	--ADDI R0,R16, x"001F"      -- INSTR 154 -- -- 
"00000000","11110000","10001000","00000101",	--AND R7,R16,R17            -- INSTR 155 -- -- LAST 5 BITS OF R7
"00000110","00010000","00000000","00000001",	--ADDI R16,R16, x"0001"     -- INSTR 156 -- -- R16 = 32 IN DECIMAL
"00000010","00010001","10001000","00000011",	--SUB R16,R17,R17           -- INSTR 157 -- -- R17 = 32 - LAST 5 BITS OF R7 
"00000010","01110011","10011000","00000011",	--SUB R19,R19,R19           -- INSTR 158 ---- ROTATION COUNTER
"00000100","00010000","00000000","00000001",	--ADDI R0,R16, x"0001"      -- INSTR 159 ---- 
"00000001","11110000","10010000","00000101",	--AND R15,R16,R18           -- INSTR 160 ---- CHECK THE LAST BIT OF R15
"00000110","01110011","00000000","00000001",	--ADDI R19,R19, x"0001"     -- INSTR 161 -- -- INCREMENT ROTATION COUNTER
"00010101","11101111","00000000","00000001",	--SHR R15,R15, x"0001"      -- INSTR 162 ---- SHIFT RIGHT BY ONE BIT
"00101010","01010000","00000000","00000010",	--BEQ R18,R16,(INSTR = 166) -- INSTR 163 -- -- IF THE LAST BIT IS 1, BRANCH TO ADDING 1 IN THE MSB
"00101010","01110001","00000000","00000100",	--BEQ R19,R17,(INSTR = 169) -- INSTR 164 --  -- END OF ROTATION CHECK
"00110000","00000000","00000000","10011111",	--JMP (INSTR = 160)         -- INSTR 165 --  -- NEXT Last bit and then SHR 
"00000001","11100011","01111000","00000001",	--ADD R15,R3,R15            -- INSTR 166 -- -- ADD x"80000000" TO R15
"00101010","01110001","00000000","00000001",	--BEQ R19,R17,(INSTR = 169) -- INSTR 167    -- END OF ROTATION CHECK
"00110000","00000000","00000000","10011111",	--JMP (INSTR = 160)         -- INSTR 168    -- NEXT SHR
"00000100","10000100","00000000","00000001",	--ADDI R4,R4, x"0001"       -- INSTR 169   -- NUMBER OF TIMES ROTATION IS CALLED
"00000000","10010000","10000000","00000101",	--AND R4,R16,R16            -- INSTR 170   -- LAST BIT OF R4
"00110000","00000000","00000000","10000110"		--JMP (INSTR = 135)         -- INSTR 171  -- JUMP BACK TO MAIN ROUTINE




);

begin

RD <= imem(CONV_INTEGER(A))&imem(CONV_INTEGER(A)+1)&imem(CONV_INTEGER(A)+2)&imem(CONV_INTEGER(A)+3);

end Behavioral;


